.title dual rc ladder
* file name rcrcac.cir
*R1 int in 10k
*V1 in 0 dc 0 ac 1 PULSE (0 5 1u 1u 1u 1 1)
*R2 out int 1k
*C1 int 0 1u
*C2 out 0 100n

Q3 A B C BJTNAME 1.0
Q4 A B C D BJTNAME 2.0
Q5 A B C D E BJTNAME 3.0

.MODEL BJTNAME NPN(BF=200 CJC=20pf CJE=20pf IS=1E-16)

.plot dc 1 2 3 4 5 6 7 8

*.control
*ac dec 10 1 100k
*plot vdb(out)
*plot ph(out)
*.endc


